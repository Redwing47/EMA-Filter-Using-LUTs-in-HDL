module ema_lut_beta (
    input  wire [7:0] addr,
    output reg  [15:0] data
);

    always @(*) begin
        case (addr)
            8'd0: data = 16'd0;
            8'd1: data = 16'd0;
            8'd2: data = 16'd1;
            8'd3: data = 16'd2;
            8'd4: data = 16'd3;
            8'd5: data = 16'd3;
            8'd6: data = 16'd4;
            8'd7: data = 16'd5;
            8'd8: data = 16'd6;
            8'd9: data = 16'd6;
            8'd10: data = 16'd7;
            8'd11: data = 16'd8;
            8'd12: data = 16'd9;
            8'd13: data = 16'd9;
            8'd14: data = 16'd10;
            8'd15: data = 16'd11;
            8'd16: data = 16'd12;
            8'd17: data = 16'd12;
            8'd18: data = 16'd13;
            8'd19: data = 16'd14;
            8'd20: data = 16'd15;
            8'd21: data = 16'd15;
            8'd22: data = 16'd16;
            8'd23: data = 16'd17;
            8'd24: data = 16'd18;
            8'd25: data = 16'd18;
            8'd26: data = 16'd19;
            8'd27: data = 16'd20;
            8'd28: data = 16'd21;
            8'd29: data = 16'd21;
            8'd30: data = 16'd22;
            8'd31: data = 16'd23;
            8'd32: data = 16'd24;
            8'd33: data = 16'd24;
            8'd34: data = 16'd25;
            8'd35: data = 16'd26;
            8'd36: data = 16'd27;
            8'd37: data = 16'd27;
            8'd38: data = 16'd28;
            8'd39: data = 16'd29;
            8'd40: data = 16'd30;
            8'd41: data = 16'd30;
            8'd42: data = 16'd31;
            8'd43: data = 16'd32;
            8'd44: data = 16'd33;
            8'd45: data = 16'd33;
            8'd46: data = 16'd34;
            8'd47: data = 16'd35;
            8'd48: data = 16'd36;
            8'd49: data = 16'd36;
            8'd50: data = 16'd37;
            8'd51: data = 16'd38;
            8'd52: data = 16'd39;
            8'd53: data = 16'd39;
            8'd54: data = 16'd40;
            8'd55: data = 16'd41;
            8'd56: data = 16'd42;
            8'd57: data = 16'd42;
            8'd58: data = 16'd43;
            8'd59: data = 16'd44;
            8'd60: data = 16'd45;
            8'd61: data = 16'd45;
            8'd62: data = 16'd46;
            8'd63: data = 16'd47;
            8'd64: data = 16'd48;
            8'd65: data = 16'd48;
            8'd66: data = 16'd49;
            8'd67: data = 16'd50;
            8'd68: data = 16'd51;
            8'd69: data = 16'd51;
            8'd70: data = 16'd52;
            8'd71: data = 16'd53;
            8'd72: data = 16'd54;
            8'd73: data = 16'd54;
            8'd74: data = 16'd55;
            8'd75: data = 16'd56;
            8'd76: data = 16'd57;
            8'd77: data = 16'd57;
            8'd78: data = 16'd58;
            8'd79: data = 16'd59;
            8'd80: data = 16'd60;
            8'd81: data = 16'd60;
            8'd82: data = 16'd61;
            8'd83: data = 16'd62;
            8'd84: data = 16'd63;
            8'd85: data = 16'd63;
            8'd86: data = 16'd64;
            8'd87: data = 16'd65;
            8'd88: data = 16'd66;
            8'd89: data = 16'd66;
            8'd90: data = 16'd67;
            8'd91: data = 16'd68;
            8'd92: data = 16'd69;
            8'd93: data = 16'd69;
            8'd94: data = 16'd70;
            8'd95: data = 16'd71;
            8'd96: data = 16'd72;
            8'd97: data = 16'd72;
            8'd98: data = 16'd73;
            8'd99: data = 16'd74;
            8'd100: data = 16'd75;
            8'd101: data = 16'd75;
            8'd102: data = 16'd76;
            8'd103: data = 16'd77;
            8'd104: data = 16'd78;
            8'd105: data = 16'd78;
            8'd106: data = 16'd79;
            8'd107: data = 16'd80;
            8'd108: data = 16'd81;
            8'd109: data = 16'd81;
            8'd110: data = 16'd82;
            8'd111: data = 16'd83;
            8'd112: data = 16'd84;
            8'd113: data = 16'd84;
            8'd114: data = 16'd85;
            8'd115: data = 16'd86;
            8'd116: data = 16'd87;
            8'd117: data = 16'd87;
            8'd118: data = 16'd88;
            8'd119: data = 16'd89;
            8'd120: data = 16'd90;
            8'd121: data = 16'd90;
            8'd122: data = 16'd91;
            8'd123: data = 16'd92;
            8'd124: data = 16'd93;
            8'd125: data = 16'd93;
            8'd126: data = 16'd94;
            8'd127: data = 16'd95;
            8'd128: data = 16'd96;
            8'd129: data = 16'd96;
            8'd130: data = 16'd97;
            8'd131: data = 16'd98;
            8'd132: data = 16'd99;
            8'd133: data = 16'd99;
            8'd134: data = 16'd100;
            8'd135: data = 16'd101;
            8'd136: data = 16'd102;
            8'd137: data = 16'd102;
            8'd138: data = 16'd103;
            8'd139: data = 16'd104;
            8'd140: data = 16'd105;
            8'd141: data = 16'd105;
            8'd142: data = 16'd106;
            8'd143: data = 16'd107;
            8'd144: data = 16'd108;
            8'd145: data = 16'd108;
            8'd146: data = 16'd109;
            8'd147: data = 16'd110;
            8'd148: data = 16'd111;
            8'd149: data = 16'd111;
            8'd150: data = 16'd112;
            8'd151: data = 16'd113;
            8'd152: data = 16'd114;
            8'd153: data = 16'd114;
            8'd154: data = 16'd115;
            8'd155: data = 16'd116;
            8'd156: data = 16'd117;
            8'd157: data = 16'd117;
            8'd158: data = 16'd118;
            8'd159: data = 16'd119;
            8'd160: data = 16'd120;
            8'd161: data = 16'd120;
            8'd162: data = 16'd121;
            8'd163: data = 16'd122;
            8'd164: data = 16'd123;
            8'd165: data = 16'd123;
            8'd166: data = 16'd124;
            8'd167: data = 16'd125;
            8'd168: data = 16'd126;
            8'd169: data = 16'd126;
            8'd170: data = 16'd127;
            8'd171: data = 16'd128;
            8'd172: data = 16'd129;
            8'd173: data = 16'd129;
            8'd174: data = 16'd130;
            8'd175: data = 16'd131;
            8'd176: data = 16'd132;
            8'd177: data = 16'd132;
            8'd178: data = 16'd133;
            8'd179: data = 16'd134;
            8'd180: data = 16'd135;
            8'd181: data = 16'd135;
            8'd182: data = 16'd136;
            8'd183: data = 16'd137;
            8'd184: data = 16'd138;
            8'd185: data = 16'd138;
            8'd186: data = 16'd139;
            8'd187: data = 16'd140;
            8'd188: data = 16'd141;
            8'd189: data = 16'd141;
            8'd190: data = 16'd142;
            8'd191: data = 16'd143;
            8'd192: data = 16'd144;
            8'd193: data = 16'd144;
            8'd194: data = 16'd145;
            8'd195: data = 16'd146;
            8'd196: data = 16'd147;
            8'd197: data = 16'd147;
            8'd198: data = 16'd148;
            8'd199: data = 16'd149;
            8'd200: data = 16'd150;
            8'd201: data = 16'd150;
            8'd202: data = 16'd151;
            8'd203: data = 16'd152;
            8'd204: data = 16'd153;
            8'd205: data = 16'd153;
            8'd206: data = 16'd154;
            8'd207: data = 16'd155;
            8'd208: data = 16'd156;
            8'd209: data = 16'd156;
            8'd210: data = 16'd157;
            8'd211: data = 16'd158;
            8'd212: data = 16'd159;
            8'd213: data = 16'd159;
            8'd214: data = 16'd160;
            8'd215: data = 16'd161;
            8'd216: data = 16'd162;
            8'd217: data = 16'd162;
            8'd218: data = 16'd163;
            8'd219: data = 16'd164;
            8'd220: data = 16'd165;
            8'd221: data = 16'd165;
            8'd222: data = 16'd166;
            8'd223: data = 16'd167;
            8'd224: data = 16'd168;
            8'd225: data = 16'd168;
            8'd226: data = 16'd169;
            8'd227: data = 16'd170;
            8'd228: data = 16'd171;
            8'd229: data = 16'd171;
            8'd230: data = 16'd172;
            8'd231: data = 16'd173;
            8'd232: data = 16'd174;
            8'd233: data = 16'd174;
            8'd234: data = 16'd175;
            8'd235: data = 16'd176;
            8'd236: data = 16'd177;
            8'd237: data = 16'd177;
            8'd238: data = 16'd178;
            8'd239: data = 16'd179;
            8'd240: data = 16'd180;
            8'd241: data = 16'd180;
            8'd242: data = 16'd181;
            8'd243: data = 16'd182;
            8'd244: data = 16'd183;
            8'd245: data = 16'd183;
            8'd246: data = 16'd184;
            8'd247: data = 16'd185;
            8'd248: data = 16'd186;
            8'd249: data = 16'd186;
            8'd250: data = 16'd187;
            8'd251: data = 16'd188;
            8'd252: data = 16'd189;
            8'd253: data = 16'd189;
            8'd254: data = 16'd190;
            8'd255: data = 16'd191;
        endcase
    end

endmodule
